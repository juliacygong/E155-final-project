// sharp symbol 
// 10 x 16

module sharp_rom (
    input logic clk,
    input logic [7:0] addr,
    output logic pixel_out
);


endmodule