// D5# LUT
// 11/5/2025
// LUT for D5# sin signal, used in simulation

module dfiveshLUT (
    input logic [8:0] add_rd,
    output logic [15:0] din
);

    (* rom_style = "distributed" *)   // For Lattice LSE
    logic [15:0] din_out;

    assign din = din_out;
    // Using a combinatorial case statement forces the synthesizer
    // to implement this as Distributed Logic (LUTs) rather than Block RAM.
    // This results in ZERO read latency.
    always_comb begin
        case (add_rd)
            9'd0: din_out = 16'b0000000010000000; //80
            9'd1: din_out = 16'b0000000011011001; //d9
            9'd2: din_out = 16'b0000000011111111; //ff
            9'd3: din_out = 16'b0000000011011011; //db
            9'd4: din_out = 16'b0000000010000011; //83
            9'd5: din_out = 16'b0000000000101001; //29
            9'd6: din_out = 16'b0000000000000001;
            9'd7: din_out = 16'b0000000000100010;
            9'd8: din_out = 16'b0000000001111010;
            9'd9: din_out = 16'b0000000011010101;
            9'd10: din_out = 16'b0000000011111111;
            9'd11: din_out = 16'b0000000011100000;
            9'd12: din_out = 16'b0000000010001010;
            9'd13: din_out = 16'b0000000000101110;
            9'd14: din_out = 16'b0000000000000001;
            9'd15: din_out = 16'b0000000000011110;
            9'd16: din_out = 16'b0000000001110011;
            9'd17: din_out = 16'b0000000011010000;
            9'd18: din_out = 16'b0000000011111110;
            9'd19: din_out = 16'b0000000011100100;
            9'd20: din_out = 16'b0000000010010000;
            9'd21: din_out = 16'b0000000000110011;
            9'd22: din_out = 16'b0000000000000010;
            9'd23: din_out = 16'b0000000000011010;
            9'd24: din_out = 16'b0000000001101101;
            9'd25: din_out = 16'b0000000011001011;
            9'd26: din_out = 16'b0000000011111101;
            9'd27: din_out = 16'b0000000011101000;
            9'd28: din_out = 16'b0000000010010110;
            9'd29: din_out = 16'b0000000000111000;
            9'd30: din_out = 16'b0000000000000011;
            9'd31: din_out = 16'b0000000000010111;
            9'd32: din_out = 16'b0000000001100111;
            9'd33: din_out = 16'b0000000011000101;
            9'd34: din_out = 16'b0000000011111100;
            9'd35: din_out = 16'b0000000011101011;
            9'd36: din_out = 16'b0000000010011100;
            9'd37: din_out = 16'b0000000000111101;
            9'd38: din_out = 16'b0000000000000101;
            9'd39: din_out = 16'b0000000000010011;
            9'd40: din_out = 16'b0000000001100000;
            9'd41: din_out = 16'b0000000011000000;
            9'd42: din_out = 16'b0000000011111011;
            9'd43: din_out = 16'b0000000011101111;
            9'd44: din_out = 16'b0000000010100011;
            9'd45: din_out = 16'b0000000001000011;
            9'd46: din_out = 16'b0000000000000110;
            9'd47: din_out = 16'b0000000000010000;
            9'd48: din_out = 16'b0000000001011010;
            9'd49: din_out = 16'b0000000010111010;
            9'd50: din_out = 16'b0000000011111001;
            9'd51: din_out = 16'b0000000011110010;
            9'd52: din_out = 16'b0000000010101001;
            9'd53: din_out = 16'b0000000001001000;
            9'd54: din_out = 16'b0000000000001000;
            9'd55: din_out = 16'b0000000000001101;
            9'd56: din_out = 16'b0000000001010100;
            9'd57: din_out = 16'b0000000010110101;
            9'd58: din_out = 16'b0000000011110111;
            9'd59: din_out = 16'b0000000011110100;
            9'd60: din_out = 16'b0000000010101111;
            9'd61: din_out = 16'b0000000001001110;
            9'd62: din_out = 16'b0000000000001011;
            9'd63: din_out = 16'b0000000000001011;
            9'd64: din_out = 16'b0000000001001110;
            9'd65: din_out = 16'b0000000010101111;
            9'd66: din_out = 16'b0000000011110100;
            9'd67: din_out = 16'b0000000011110111;
            9'd68: din_out = 16'b0000000010110101;
            9'd69: din_out = 16'b0000000001010100;
            9'd70: din_out = 16'b0000000000001101;
            9'd71: din_out = 16'b0000000000001000;
            9'd72: din_out = 16'b0000000001001000;
            9'd73: din_out = 16'b0000000010101001;
            9'd74: din_out = 16'b0000000011110010;
            9'd75: din_out = 16'b0000000011111001;
            9'd76: din_out = 16'b0000000010111010;
            9'd77: din_out = 16'b0000000001011010;
            9'd78: din_out = 16'b0000000000010000;
            9'd79: din_out = 16'b0000000000000110;
            9'd80: din_out = 16'b0000000001000011;
            9'd81: din_out = 16'b0000000010100011;
            9'd82: din_out = 16'b0000000011101111;
            9'd83: din_out = 16'b0000000011111011;
            9'd84: din_out = 16'b0000000011000000;
            9'd85: din_out = 16'b0000000001100000;
            9'd86: din_out = 16'b0000000000010011;
            9'd87: din_out = 16'b0000000000000101;
            9'd88: din_out = 16'b0000000000111101;
            9'd89: din_out = 16'b0000000010011100;
            9'd90: din_out = 16'b0000000011101011;
            9'd91: din_out = 16'b0000000011111100;
            9'd92: din_out = 16'b0000000011000101;
            9'd93: din_out = 16'b0000000001100111;
            9'd94: din_out = 16'b0000000000010111;
            9'd95: din_out = 16'b0000000000000011;
            9'd96: din_out = 16'b0000000000111000;
            9'd97: din_out = 16'b0000000010010110;
            9'd98: din_out = 16'b0000000011101000;
            9'd99: din_out = 16'b0000000011111101;
            9'd100: din_out = 16'b0000000011001011;
            9'd101: din_out = 16'b0000000001101101;
            9'd102: din_out = 16'b0000000000011010;
            9'd103: din_out = 16'b0000000000000010;
            9'd104: din_out = 16'b0000000000110011;
            9'd105: din_out = 16'b0000000010010000;
            9'd106: din_out = 16'b0000000011100100;
            9'd107: din_out = 16'b0000000011111110;
            9'd108: din_out = 16'b0000000011010000;
            9'd109: din_out = 16'b0000000001110011;
            9'd110: din_out = 16'b0000000000011110;
            9'd111: din_out = 16'b0000000000000001;
            9'd112: din_out = 16'b0000000000101110;
            9'd113: din_out = 16'b0000000010001010;
            9'd114: din_out = 16'b0000000011100000;
            9'd115: din_out = 16'b0000000011111111;
            9'd116: din_out = 16'b0000000011010101;
            9'd117: din_out = 16'b0000000001111010;
            9'd118: din_out = 16'b0000000000100010;
            9'd119: din_out = 16'b0000000000000001;
            9'd120: din_out = 16'b0000000000101001;
            9'd121: din_out = 16'b0000000010000011;
            9'd122: din_out = 16'b0000000011011011;
            9'd123: din_out = 16'b0000000011111111;
            9'd124: din_out = 16'b0000000011011001;
            9'd125: din_out = 16'b0000000010000000;
            9'd126: din_out = 16'b0000000000100111;
            9'd127: din_out = 16'b0000000000000001;
            9'd128: din_out = 16'b0000000000100101;
            9'd129: din_out = 16'b0000000001111101;
            9'd130: din_out = 16'b0000000011010111;
            9'd131: din_out = 16'b0000000011111111;
            9'd132: din_out = 16'b0000000011011110;
            9'd133: din_out = 16'b0000000010000110;
            9'd134: din_out = 16'b0000000000101011;
            9'd135: din_out = 16'b0000000000000001;
            9'd136: din_out = 16'b0000000000100000;
            9'd137: din_out = 16'b0000000001110110;
            9'd138: din_out = 16'b0000000011010010;
            9'd139: din_out = 16'b0000000011111111;
            9'd140: din_out = 16'b0000000011100010;
            9'd141: din_out = 16'b0000000010001101;
            9'd142: din_out = 16'b0000000000110000;
            9'd143: din_out = 16'b0000000000000010;
            9'd144: din_out = 16'b0000000000011100;
            9'd145: din_out = 16'b0000000001110000;
            9'd146: din_out = 16'b0000000011001101;
            9'd147: din_out = 16'b0000000011111110;
            9'd148: din_out = 16'b0000000011100110;
            9'd149: din_out = 16'b0000000010010011;
            9'd150: din_out = 16'b0000000000110101;
            9'd151: din_out = 16'b0000000000000011;
            9'd152: din_out = 16'b0000000000011000;
            9'd153: din_out = 16'b0000000001101010;
            9'd154: din_out = 16'b0000000011001000;
            9'd155: din_out = 16'b0000000011111101;
            9'd156: din_out = 16'b0000000011101001;
            9'd157: din_out = 16'b0000000010011001;
            9'd158: din_out = 16'b0000000000111011;
            9'd159: din_out = 16'b0000000000000100;
            9'd160: din_out = 16'b0000000000010101;
            9'd161: din_out = 16'b0000000001100100;
            9'd162: din_out = 16'b0000000011000011;
            9'd163: din_out = 16'b0000000011111011;
            9'd164: din_out = 16'b0000000011101101;
            9'd165: din_out = 16'b0000000010100000;
            9'd166: din_out = 16'b0000000001000000;
            9'd167: din_out = 16'b0000000000000101;
            9'd168: din_out = 16'b0000000000010001;
            9'd169: din_out = 16'b0000000001011101;
            9'd170: din_out = 16'b0000000010111101;
            9'd171: din_out = 16'b0000000011111010;
            9'd172: din_out = 16'b0000000011110000;
            9'd173: din_out = 16'b0000000010100110;
            9'd174: din_out = 16'b0000000001000110;
            9'd175: din_out = 16'b0000000000000111;
            9'd176: din_out = 16'b0000000000001110;
            9'd177: din_out = 16'b0000000001010111;
            9'd178: din_out = 16'b0000000010111000;
            9'd179: din_out = 16'b0000000011111000;
            9'd180: din_out = 16'b0000000011110011;
            9'd181: din_out = 16'b0000000010101100;
            9'd182: din_out = 16'b0000000001001011;
            9'd183: din_out = 16'b0000000000001001;
            9'd184: din_out = 16'b0000000000001100;
            9'd185: din_out = 16'b0000000001010001;
            9'd186: din_out = 16'b0000000010110010;
            9'd187: din_out = 16'b0000000011110101;
            9'd188: din_out = 16'b0000000011110101;
            9'd189: din_out = 16'b0000000010110010;
            9'd190: din_out = 16'b0000000001010001;
            9'd191: din_out = 16'b0000000000001100;
            9'd192: din_out = 16'b0000000000001001;
            9'd193: din_out = 16'b0000000001001011;
            9'd194: din_out = 16'b0000000010101100;
            9'd195: din_out = 16'b0000000011110011;
            9'd196: din_out = 16'b0000000011111000;
            9'd197: din_out = 16'b0000000010111000;
            9'd198: din_out = 16'b0000000001010111;
            9'd199: din_out = 16'b0000000000001110;
            9'd200: din_out = 16'b0000000000000111;
            9'd201: din_out = 16'b0000000001000110;
            9'd202: din_out = 16'b0000000010100110;
            9'd203: din_out = 16'b0000000011110000;
            9'd204: din_out = 16'b0000000011111010;
            9'd205: din_out = 16'b0000000010111101;
            9'd206: din_out = 16'b0000000001011101;
            9'd207: din_out = 16'b0000000000010001;
            9'd208: din_out = 16'b0000000000000101;
            9'd209: din_out = 16'b0000000001000000;
            9'd210: din_out = 16'b0000000010100000;
            9'd211: din_out = 16'b0000000011101101;
            9'd212: din_out = 16'b0000000011111011;
            9'd213: din_out = 16'b0000000011000011;
            9'd214: din_out = 16'b0000000001100100;
            9'd215: din_out = 16'b0000000000010101;
            9'd216: din_out = 16'b0000000000000100;
            9'd217: din_out = 16'b0000000000111011;
            9'd218: din_out = 16'b0000000010011001;
            9'd219: din_out = 16'b0000000011101001;
            9'd220: din_out = 16'b0000000011111101;
            9'd221: din_out = 16'b0000000011001000;
            9'd222: din_out = 16'b0000000001101010;
            9'd223: din_out = 16'b0000000000011000;
            9'd224: din_out = 16'b0000000000000011;
            9'd225: din_out = 16'b0000000000110101;
            9'd226: din_out = 16'b0000000010010011;
            9'd227: din_out = 16'b0000000011100110;
            9'd228: din_out = 16'b0000000011111110;
            9'd229: din_out = 16'b0000000011001101;
            9'd230: din_out = 16'b0000000001110000;
            9'd231: din_out = 16'b0000000000011100;
            9'd232: din_out = 16'b0000000000000010;
            9'd233: din_out = 16'b0000000000110000;
            9'd234: din_out = 16'b0000000010001101;
            9'd235: din_out = 16'b0000000011100010;
            9'd236: din_out = 16'b0000000011111111;
            9'd237: din_out = 16'b0000000011010010;
            9'd238: din_out = 16'b0000000001110110;
            9'd239: din_out = 16'b0000000000100000;
            9'd240: din_out = 16'b0000000000000001;
            9'd241: din_out = 16'b0000000000101011;
            9'd242: din_out = 16'b0000000010000110;
            9'd243: din_out = 16'b0000000011011110;
            9'd244: din_out = 16'b0000000011111111;
            9'd245: din_out = 16'b0000000011010111;
            9'd246: din_out = 16'b0000000001111101;
            9'd247: din_out = 16'b0000000000100101;
            9'd248: din_out = 16'b0000000000000001;
            9'd249: din_out = 16'b0000000000100111;
            9'd250: din_out = 16'b0000000010000000;
            9'd251: din_out = 16'b0000000011011001;
            9'd252: din_out = 16'b0000000011111111;
            9'd253: din_out = 16'b0000000011011011;
            9'd254: din_out = 16'b0000000010000011;
            9'd255: din_out = 16'b0000000000101001;
            9'd256: din_out = 16'b0000000000000001;
            9'd257: din_out = 16'b0000000000100010;
            9'd258: din_out = 16'b0000000001111010;
            9'd259: din_out = 16'b0000000011010101;
            9'd260: din_out = 16'b0000000011111111;
            9'd261: din_out = 16'b0000000011100000;
            9'd262: din_out = 16'b0000000010001010;
            9'd263: din_out = 16'b0000000000101110;
            9'd264: din_out = 16'b0000000000000001;
            9'd265: din_out = 16'b0000000000011110;
            9'd266: din_out = 16'b0000000001110011;
            9'd267: din_out = 16'b0000000011010000;
            9'd268: din_out = 16'b0000000011111110;
            9'd269: din_out = 16'b0000000011100100;
            9'd270: din_out = 16'b0000000010010000;
            9'd271: din_out = 16'b0000000000110011;
            9'd272: din_out = 16'b0000000000000010;
            9'd273: din_out = 16'b0000000000011010;
            9'd274: din_out = 16'b0000000001101101;
            9'd275: din_out = 16'b0000000011001011;
            9'd276: din_out = 16'b0000000011111101;
            9'd277: din_out = 16'b0000000011101000;
            9'd278: din_out = 16'b0000000010010110;
            9'd279: din_out = 16'b0000000000111000;
            9'd280: din_out = 16'b0000000000000011;
            9'd281: din_out = 16'b0000000000010111;
            9'd282: din_out = 16'b0000000001100111;
            9'd283: din_out = 16'b0000000011000101;
            9'd284: din_out = 16'b0000000011111100;
            9'd285: din_out = 16'b0000000011101011;
            9'd286: din_out = 16'b0000000010011100;
            9'd287: din_out = 16'b0000000000111101;
            9'd288: din_out = 16'b0000000000000101;
            9'd289: din_out = 16'b0000000000010011;
            9'd290: din_out = 16'b0000000001100000;
            9'd291: din_out = 16'b0000000011000000;
            9'd292: din_out = 16'b0000000011111011;
            9'd293: din_out = 16'b0000000011101111;
            9'd294: din_out = 16'b0000000010100011;
            9'd295: din_out = 16'b0000000001000011;
            9'd296: din_out = 16'b0000000000000110;
            9'd297: din_out = 16'b0000000000010000;
            9'd298: din_out = 16'b0000000001011010;
            9'd299: din_out = 16'b0000000010111010;
            9'd300: din_out = 16'b0000000011111001;
            9'd301: din_out = 16'b0000000011110010;
            9'd302: din_out = 16'b0000000010101001;
            9'd303: din_out = 16'b0000000001001000;
            9'd304: din_out = 16'b0000000000001000;
            9'd305: din_out = 16'b0000000000001101;
            9'd306: din_out = 16'b0000000001010100;
            9'd307: din_out = 16'b0000000010110101;
            9'd308: din_out = 16'b0000000011110111;
            9'd309: din_out = 16'b0000000011110100;
            9'd310: din_out = 16'b0000000010101111;
            9'd311: din_out = 16'b0000000001001110;
            9'd312: din_out = 16'b0000000000001011;
            9'd313: din_out = 16'b0000000000001011;
            9'd314: din_out = 16'b0000000001001110;
            9'd315: din_out = 16'b0000000010101111;
            9'd316: din_out = 16'b0000000011110100;
            9'd317: din_out = 16'b0000000011110111;
            9'd318: din_out = 16'b0000000010110101;
            9'd319: din_out = 16'b0000000001010100;
            9'd320: din_out = 16'b0000000000001101;
            9'd321: din_out = 16'b0000000000001000;
            9'd322: din_out = 16'b0000000001001000;
            9'd323: din_out = 16'b0000000010101001;
            9'd324: din_out = 16'b0000000011110010;
            9'd325: din_out = 16'b0000000011111001;
            9'd326: din_out = 16'b0000000010111010;
            9'd327: din_out = 16'b0000000001011010;
            9'd328: din_out = 16'b0000000000010000;
            9'd329: din_out = 16'b0000000000000110;
            9'd330: din_out = 16'b0000000001000011;
            9'd331: din_out = 16'b0000000010100011;
            9'd332: din_out = 16'b0000000011101111;
            9'd333: din_out = 16'b0000000011111011;
            9'd334: din_out = 16'b0000000011000000;
            9'd335: din_out = 16'b0000000001100000;
            9'd336: din_out = 16'b0000000000010011;
            9'd337: din_out = 16'b0000000000000101;
            9'd338: din_out = 16'b0000000000111101;
            9'd339: din_out = 16'b0000000010011100;
            9'd340: din_out = 16'b0000000011101011;
            9'd341: din_out = 16'b0000000011111100;
            9'd342: din_out = 16'b0000000011000101;
            9'd343: din_out = 16'b0000000001100111;
            9'd344: din_out = 16'b0000000000010111;
            9'd345: din_out = 16'b0000000000000011;
            9'd346: din_out = 16'b0000000000111000;
            9'd347: din_out = 16'b0000000010010110;
            9'd348: din_out = 16'b0000000011101000;
            9'd349: din_out = 16'b0000000011111101;
            9'd350: din_out = 16'b0000000011001011;
            9'd351: din_out = 16'b0000000001101101;
            9'd352: din_out = 16'b0000000000011010;
            9'd353: din_out = 16'b0000000000000010;
            9'd354: din_out = 16'b0000000000110011;
            9'd355: din_out = 16'b0000000010010000;
            9'd356: din_out = 16'b0000000011100100;
            9'd357: din_out = 16'b0000000011111110;
            9'd358: din_out = 16'b0000000011010000;
            9'd359: din_out = 16'b0000000001110011;
            9'd360: din_out = 16'b0000000000011110;
            9'd361: din_out = 16'b0000000000000001;
            9'd362: din_out = 16'b0000000000101110;
            9'd363: din_out = 16'b0000000010001010;
            9'd364: din_out = 16'b0000000011100000;
            9'd365: din_out = 16'b0000000011111111;
            9'd366: din_out = 16'b0000000011010101;
            9'd367: din_out = 16'b0000000001111010;
            9'd368: din_out = 16'b0000000000100010;
            9'd369: din_out = 16'b0000000000000001;
            9'd370: din_out = 16'b0000000000101001;
            9'd371: din_out = 16'b0000000010000011;
            9'd372: din_out = 16'b0000000011011011;
            9'd373: din_out = 16'b0000000011111111;
            9'd374: din_out = 16'b0000000011011001;
            9'd375: din_out = 16'b0000000010000000;
            9'd376: din_out = 16'b0000000000100111;
            9'd377: din_out = 16'b0000000000000001;
            9'd378: din_out = 16'b0000000000100101;
            9'd379: din_out = 16'b0000000001111101;
            9'd380: din_out = 16'b0000000011010111;
            9'd381: din_out = 16'b0000000011111111;
            9'd382: din_out = 16'b0000000011011110;
            9'd383: din_out = 16'b0000000010000110;
            9'd384: din_out = 16'b0000000000101011;
            9'd385: din_out = 16'b0000000000000001;
            9'd386: din_out = 16'b0000000000100000;
            9'd387: din_out = 16'b0000000001110110;
            9'd388: din_out = 16'b0000000011010010;
            9'd389: din_out = 16'b0000000011111111;
            9'd390: din_out = 16'b0000000011100010;
            9'd391: din_out = 16'b0000000010001101;
            9'd392: din_out = 16'b0000000000110000;
            9'd393: din_out = 16'b0000000000000010;
            9'd394: din_out = 16'b0000000000011100;
            9'd395: din_out = 16'b0000000001110000;
            9'd396: din_out = 16'b0000000011001101;
            9'd397: din_out = 16'b0000000011111110;
            9'd398: din_out = 16'b0000000011100110;
            9'd399: din_out = 16'b0000000010010011;
            9'd400: din_out = 16'b0000000000110101;
            9'd401: din_out = 16'b0000000000000011;
            9'd402: din_out = 16'b0000000000011000;
            9'd403: din_out = 16'b0000000001101010;
            9'd404: din_out = 16'b0000000011001000;
            9'd405: din_out = 16'b0000000011111101;
            9'd406: din_out = 16'b0000000011101001;
            9'd407: din_out = 16'b0000000010011001;
            9'd408: din_out = 16'b0000000000111011;
            9'd409: din_out = 16'b0000000000000100;
            9'd410: din_out = 16'b0000000000010101;
            9'd411: din_out = 16'b0000000001100100;
            9'd412: din_out = 16'b0000000011000011;
            9'd413: din_out = 16'b0000000011111011;
            9'd414: din_out = 16'b0000000011101101;
            9'd415: din_out = 16'b0000000010100000;
            9'd416: din_out = 16'b0000000001000000;
            9'd417: din_out = 16'b0000000000000101;
            9'd418: din_out = 16'b0000000000010001;
            9'd419: din_out = 16'b0000000001011101;
            9'd420: din_out = 16'b0000000010111101;
            9'd421: din_out = 16'b0000000011111010;
            9'd422: din_out = 16'b0000000011110000;
            9'd423: din_out = 16'b0000000010100110;
            9'd424: din_out = 16'b0000000001000110;
            9'd425: din_out = 16'b0000000000000111;
            9'd426: din_out = 16'b0000000000001110;
            9'd427: din_out = 16'b0000000001010111;
            9'd428: din_out = 16'b0000000010111000;
            9'd429: din_out = 16'b0000000011111000;
            9'd430: din_out = 16'b0000000011110011;
            9'd431: din_out = 16'b0000000010101100;
            9'd432: din_out = 16'b0000000001001011;
            9'd433: din_out = 16'b0000000000001001;
            9'd434: din_out = 16'b0000000000001100;
            9'd435: din_out = 16'b0000000001010001;
            9'd436: din_out = 16'b0000000010110010;
            9'd437: din_out = 16'b0000000011110101;
            9'd438: din_out = 16'b0000000011110101;
            9'd439: din_out = 16'b0000000010110010;
            9'd440: din_out = 16'b0000000001010001;
            9'd441: din_out = 16'b0000000000001100;
            9'd442: din_out = 16'b0000000000001001;
            9'd443: din_out = 16'b0000000001001011;
            9'd444: din_out = 16'b0000000010101100;
            9'd445: din_out = 16'b0000000011110011;
            9'd446: din_out = 16'b0000000011111000;
            9'd447: din_out = 16'b0000000010111000;
            9'd448: din_out = 16'b0000000001010111;
            9'd449: din_out = 16'b0000000000001110;
            9'd450: din_out = 16'b0000000000000111;
            9'd451: din_out = 16'b0000000001000110;
            9'd452: din_out = 16'b0000000010100110;
            9'd453: din_out = 16'b0000000011110000;
            9'd454: din_out = 16'b0000000011111010;
            9'd455: din_out = 16'b0000000010111101;
            9'd456: din_out = 16'b0000000001011101;
            9'd457: din_out = 16'b0000000000010001;
            9'd458: din_out = 16'b0000000000000101;
            9'd459: din_out = 16'b0000000001000000;
            9'd460: din_out = 16'b0000000010100000;
            9'd461: din_out = 16'b0000000011101101;
            9'd462: din_out = 16'b0000000011111011;
            9'd463: din_out = 16'b0000000011000011;
            9'd464: din_out = 16'b0000000001100100;
            9'd465: din_out = 16'b0000000000010101;
            9'd466: din_out = 16'b0000000000000100;
            9'd467: din_out = 16'b0000000000111011;
            9'd468: din_out = 16'b0000000010011001;
            9'd469: din_out = 16'b0000000011101001;
            9'd470: din_out = 16'b0000000011111101;
            9'd471: din_out = 16'b0000000011001000;
            9'd472: din_out = 16'b0000000001101010;
            9'd473: din_out = 16'b0000000000011000;
            9'd474: din_out = 16'b0000000000000011;
            9'd475: din_out = 16'b0000000000110101;
            9'd476: din_out = 16'b0000000010010011;
            9'd477: din_out = 16'b0000000011100110;
            9'd478: din_out = 16'b0000000011111110;
            9'd479: din_out = 16'b0000000011001101;
            9'd480: din_out = 16'b0000000001110000;
            9'd481: din_out = 16'b0000000000011100;
            9'd482: din_out = 16'b0000000000000010;
            9'd483: din_out = 16'b0000000000110000;
            9'd484: din_out = 16'b0000000010001101;
            9'd485: din_out = 16'b0000000011100010;
            9'd486: din_out = 16'b0000000011111111;
            9'd487: din_out = 16'b0000000011010010;
            9'd488: din_out = 16'b0000000001110110;
            9'd489: din_out = 16'b0000000000100000;
            9'd490: din_out = 16'b0000000000000001;
            9'd491: din_out = 16'b0000000000101011;
            9'd492: din_out = 16'b0000000010000110;
            9'd493: din_out = 16'b0000000011011110;
            9'd494: din_out = 16'b0000000011111111;
            9'd495: din_out = 16'b0000000011010111;
            9'd496: din_out = 16'b0000000001111101;
            9'd497: din_out = 16'b0000000000100101;
            9'd498: din_out = 16'b0000000000000001;
            9'd499: din_out = 16'b0000000000100111;
            9'd500: din_out = 16'b0000000010000000;
            9'd501: din_out = 16'b0000000011011001;
            9'd502: din_out = 16'b0000000011111111;
            9'd503: din_out = 16'b0000000011011011;
            9'd504: din_out = 16'b0000000010000011;
            9'd505: din_out = 16'b0000000000101001;
            9'd506: din_out = 16'b0000000000000001;
            9'd507: din_out = 16'b0000000000100010;
            9'd508: din_out = 16'b0000000001111010;
            9'd509: din_out = 16'b0000000011010101;
            9'd510: din_out = 16'b0000000011111111;
            9'd511: din_out = 16'b0000000011100000;
            default: din_out = 16'd0;
        endcase
    end

endmodule