module dfiveshLUT (input logic [8:0] add_rd,
				  output logic [15:0] din_out);

logic [511:0][15:0] din;
assign din[0] = 16'b0000000010000000;
assign din[1] = 16'b0000000011011001;
assign din[2] = 16'b0000000011111111;
assign din[3] = 16'b0000000011011011;
assign din[4] = 16'b0000000010000011;
assign din[5] = 16'b0000000000101001;
assign din[6] = 16'b0000000000000001;
assign din[7] = 16'b0000000000100010;
assign din[8] = 16'b0000000001111010;
assign din[9] = 16'b0000000011010101;
assign din[10] = 16'b0000000011111111;
assign din[11] = 16'b0000000011100000;
assign din[12] = 16'b0000000010001010;
assign din[13] = 16'b0000000000101110;
assign din[14] = 16'b0000000000000001;
assign din[15] = 16'b0000000000011110;
assign din[16] = 16'b0000000001110011;
assign din[17] = 16'b0000000011010000;
assign din[18] = 16'b0000000011111110;
assign din[19] = 16'b0000000011100100;
assign din[20] = 16'b0000000010010000;
assign din[21] = 16'b0000000000110011;
assign din[22] = 16'b0000000000000010;
assign din[23] = 16'b0000000000011010;
assign din[24] = 16'b0000000001101101;
assign din[25] = 16'b0000000011001011;
assign din[26] = 16'b0000000011111101;
assign din[27] = 16'b0000000011101000;
assign din[28] = 16'b0000000010010110;
assign din[29] = 16'b0000000000111000;
assign din[30] = 16'b0000000000000011;
assign din[31] = 16'b0000000000010111;
assign din[32] = 16'b0000000001100111;
assign din[33] = 16'b0000000011000101;
assign din[34] = 16'b0000000011111100;
assign din[35] = 16'b0000000011101011;
assign din[36] = 16'b0000000010011100;
assign din[37] = 16'b0000000000111101;
assign din[38] = 16'b0000000000000101;
assign din[39] = 16'b0000000000010011;
assign din[40] = 16'b0000000001100000;
assign din[41] = 16'b0000000011000000;
assign din[42] = 16'b0000000011111011;
assign din[43] = 16'b0000000011101111;
assign din[44] = 16'b0000000010100011;
assign din[45] = 16'b0000000001000011;
assign din[46] = 16'b0000000000000110;
assign din[47] = 16'b0000000000010000;
assign din[48] = 16'b0000000001011010;
assign din[49] = 16'b0000000010111010;
assign din[50] = 16'b0000000011111001;
assign din[51] = 16'b0000000011110010;
assign din[52] = 16'b0000000010101001;
assign din[53] = 16'b0000000001001000;
assign din[54] = 16'b0000000000001000;
assign din[55] = 16'b0000000000001101;
assign din[56] = 16'b0000000001010100;
assign din[57] = 16'b0000000010110101;
assign din[58] = 16'b0000000011110111;
assign din[59] = 16'b0000000011110100;
assign din[60] = 16'b0000000010101111;
assign din[61] = 16'b0000000001001110;
assign din[62] = 16'b0000000000001011;
assign din[63] = 16'b0000000000001011;
assign din[64] = 16'b0000000001001110;
assign din[65] = 16'b0000000010101111;
assign din[66] = 16'b0000000011110100;
assign din[67] = 16'b0000000011110111;
assign din[68] = 16'b0000000010110101;
assign din[69] = 16'b0000000001010100;
assign din[70] = 16'b0000000000001101;
assign din[71] = 16'b0000000000001000;
assign din[72] = 16'b0000000001001000;
assign din[73] = 16'b0000000010101001;
assign din[74] = 16'b0000000011110010;
assign din[75] = 16'b0000000011111001;
assign din[76] = 16'b0000000010111010;
assign din[77] = 16'b0000000001011010;
assign din[78] = 16'b0000000000010000;
assign din[79] = 16'b0000000000000110;
assign din[80] = 16'b0000000001000011;
assign din[81] = 16'b0000000010100011;
assign din[82] = 16'b0000000011101111;
assign din[83] = 16'b0000000011111011;
assign din[84] = 16'b0000000011000000;
assign din[85] = 16'b0000000001100000;
assign din[86] = 16'b0000000000010011;
assign din[87] = 16'b0000000000000101;
assign din[88] = 16'b0000000000111101;
assign din[89] = 16'b0000000010011100;
assign din[90] = 16'b0000000011101011;
assign din[91] = 16'b0000000011111100;
assign din[92] = 16'b0000000011000101;
assign din[93] = 16'b0000000001100111;
assign din[94] = 16'b0000000000010111;
assign din[95] = 16'b0000000000000011;
assign din[96] = 16'b0000000000111000;
assign din[97] = 16'b0000000010010110;
assign din[98] = 16'b0000000011101000;
assign din[99] = 16'b0000000011111101;
assign din[100] = 16'b0000000011001011;
assign din[101] = 16'b0000000001101101;
assign din[102] = 16'b0000000000011010;
assign din[103] = 16'b0000000000000010;
assign din[104] = 16'b0000000000110011;
assign din[105] = 16'b0000000010010000;
assign din[106] = 16'b0000000011100100;
assign din[107] = 16'b0000000011111110;
assign din[108] = 16'b0000000011010000;
assign din[109] = 16'b0000000001110011;
assign din[110] = 16'b0000000000011110;
assign din[111] = 16'b0000000000000001;
assign din[112] = 16'b0000000000101110;
assign din[113] = 16'b0000000010001010;
assign din[114] = 16'b0000000011100000;
assign din[115] = 16'b0000000011111111;
assign din[116] = 16'b0000000011010101;
assign din[117] = 16'b0000000001111010;
assign din[118] = 16'b0000000000100010;
assign din[119] = 16'b0000000000000001;
assign din[120] = 16'b0000000000101001;
assign din[121] = 16'b0000000010000011;
assign din[122] = 16'b0000000011011011;
assign din[123] = 16'b0000000011111111;
assign din[124] = 16'b0000000011011001;
assign din[125] = 16'b0000000010000000;
assign din[126] = 16'b0000000000100111;
assign din[127] = 16'b0000000000000001;
assign din[128] = 16'b0000000000100101;
assign din[129] = 16'b0000000001111101;
assign din[130] = 16'b0000000011010111;
assign din[131] = 16'b0000000011111111;
assign din[132] = 16'b0000000011011110;
assign din[133] = 16'b0000000010000110;
assign din[134] = 16'b0000000000101011;
assign din[135] = 16'b0000000000000001;
assign din[136] = 16'b0000000000100000;
assign din[137] = 16'b0000000001110110;
assign din[138] = 16'b0000000011010010;
assign din[139] = 16'b0000000011111111;
assign din[140] = 16'b0000000011100010;
assign din[141] = 16'b0000000010001101;
assign din[142] = 16'b0000000000110000;
assign din[143] = 16'b0000000000000010;
assign din[144] = 16'b0000000000011100;
assign din[145] = 16'b0000000001110000;
assign din[146] = 16'b0000000011001101;
assign din[147] = 16'b0000000011111110;
assign din[148] = 16'b0000000011100110;
assign din[149] = 16'b0000000010010011;
assign din[150] = 16'b0000000000110101;
assign din[151] = 16'b0000000000000011;
assign din[152] = 16'b0000000000011000;
assign din[153] = 16'b0000000001101010;
assign din[154] = 16'b0000000011001000;
assign din[155] = 16'b0000000011111101;
assign din[156] = 16'b0000000011101001;
assign din[157] = 16'b0000000010011001;
assign din[158] = 16'b0000000000111011;
assign din[159] = 16'b0000000000000100;
assign din[160] = 16'b0000000000010101;
assign din[161] = 16'b0000000001100100;
assign din[162] = 16'b0000000011000011;
assign din[163] = 16'b0000000011111011;
assign din[164] = 16'b0000000011101101;
assign din[165] = 16'b0000000010100000;
assign din[166] = 16'b0000000001000000;
assign din[167] = 16'b0000000000000101;
assign din[168] = 16'b0000000000010001;
assign din[169] = 16'b0000000001011101;
assign din[170] = 16'b0000000010111101;
assign din[171] = 16'b0000000011111010;
assign din[172] = 16'b0000000011110000;
assign din[173] = 16'b0000000010100110;
assign din[174] = 16'b0000000001000110;
assign din[175] = 16'b0000000000000111;
assign din[176] = 16'b0000000000001110;
assign din[177] = 16'b0000000001010111;
assign din[178] = 16'b0000000010111000;
assign din[179] = 16'b0000000011111000;
assign din[180] = 16'b0000000011110011;
assign din[181] = 16'b0000000010101100;
assign din[182] = 16'b0000000001001011;
assign din[183] = 16'b0000000000001001;
assign din[184] = 16'b0000000000001100;
assign din[185] = 16'b0000000001010001;
assign din[186] = 16'b0000000010110010;
assign din[187] = 16'b0000000011110101;
assign din[188] = 16'b0000000011110101;
assign din[189] = 16'b0000000010110010;
assign din[190] = 16'b0000000001010001;
assign din[191] = 16'b0000000000001100;
assign din[192] = 16'b0000000000001001;
assign din[193] = 16'b0000000001001011;
assign din[194] = 16'b0000000010101100;
assign din[195] = 16'b0000000011110011;
assign din[196] = 16'b0000000011111000;
assign din[197] = 16'b0000000010111000;
assign din[198] = 16'b0000000001010111;
assign din[199] = 16'b0000000000001110;
assign din[200] = 16'b0000000000000111;
assign din[201] = 16'b0000000001000110;
assign din[202] = 16'b0000000010100110;
assign din[203] = 16'b0000000011110000;
assign din[204] = 16'b0000000011111010;
assign din[205] = 16'b0000000010111101;
assign din[206] = 16'b0000000001011101;
assign din[207] = 16'b0000000000010001;
assign din[208] = 16'b0000000000000101;
assign din[209] = 16'b0000000001000000;
assign din[210] = 16'b0000000010100000;
assign din[211] = 16'b0000000011101101;
assign din[212] = 16'b0000000011111011;
assign din[213] = 16'b0000000011000011;
assign din[214] = 16'b0000000001100100;
assign din[215] = 16'b0000000000010101;
assign din[216] = 16'b0000000000000100;
assign din[217] = 16'b0000000000111011;
assign din[218] = 16'b0000000010011001;
assign din[219] = 16'b0000000011101001;
assign din[220] = 16'b0000000011111101;
assign din[221] = 16'b0000000011001000;
assign din[222] = 16'b0000000001101010;
assign din[223] = 16'b0000000000011000;
assign din[224] = 16'b0000000000000011;
assign din[225] = 16'b0000000000110101;
assign din[226] = 16'b0000000010010011;
assign din[227] = 16'b0000000011100110;
assign din[228] = 16'b0000000011111110;
assign din[229] = 16'b0000000011001101;
assign din[230] = 16'b0000000001110000;
assign din[231] = 16'b0000000000011100;
assign din[232] = 16'b0000000000000010;
assign din[233] = 16'b0000000000110000;
assign din[234] = 16'b0000000010001101;
assign din[235] = 16'b0000000011100010;
assign din[236] = 16'b0000000011111111;
assign din[237] = 16'b0000000011010010;
assign din[238] = 16'b0000000001110110;
assign din[239] = 16'b0000000000100000;
assign din[240] = 16'b0000000000000001;
assign din[241] = 16'b0000000000101011;
assign din[242] = 16'b0000000010000110;
assign din[243] = 16'b0000000011011110;
assign din[244] = 16'b0000000011111111;
assign din[245] = 16'b0000000011010111;
assign din[246] = 16'b0000000001111101;
assign din[247] = 16'b0000000000100101;
assign din[248] = 16'b0000000000000001;
assign din[249] = 16'b0000000000100111;
assign din[250] = 16'b0000000010000000;
assign din[251] = 16'b0000000011011001;
assign din[252] = 16'b0000000011111111;
assign din[253] = 16'b0000000011011011;
assign din[254] = 16'b0000000010000011;
assign din[255] = 16'b0000000000101001;
assign din[256] = 16'b0000000000000001;
assign din[257] = 16'b0000000000100010;
assign din[258] = 16'b0000000001111010;
assign din[259] = 16'b0000000011010101;
assign din[260] = 16'b0000000011111111;
assign din[261] = 16'b0000000011100000;
assign din[262] = 16'b0000000010001010;
assign din[263] = 16'b0000000000101110;
assign din[264] = 16'b0000000000000001;
assign din[265] = 16'b0000000000011110;
assign din[266] = 16'b0000000001110011;
assign din[267] = 16'b0000000011010000;
assign din[268] = 16'b0000000011111110;
assign din[269] = 16'b0000000011100100;
assign din[270] = 16'b0000000010010000;
assign din[271] = 16'b0000000000110011;
assign din[272] = 16'b0000000000000010;
assign din[273] = 16'b0000000000011010;
assign din[274] = 16'b0000000001101101;
assign din[275] = 16'b0000000011001011;
assign din[276] = 16'b0000000011111101;
assign din[277] = 16'b0000000011101000;
assign din[278] = 16'b0000000010010110;
assign din[279] = 16'b0000000000111000;
assign din[280] = 16'b0000000000000011;
assign din[281] = 16'b0000000000010111;
assign din[282] = 16'b0000000001100111;
assign din[283] = 16'b0000000011000101;
assign din[284] = 16'b0000000011111100;
assign din[285] = 16'b0000000011101011;
assign din[286] = 16'b0000000010011100;
assign din[287] = 16'b0000000000111101;
assign din[288] = 16'b0000000000000101;
assign din[289] = 16'b0000000000010011;
assign din[290] = 16'b0000000001100000;
assign din[291] = 16'b0000000011000000;
assign din[292] = 16'b0000000011111011;
assign din[293] = 16'b0000000011101111;
assign din[294] = 16'b0000000010100011;
assign din[295] = 16'b0000000001000011;
assign din[296] = 16'b0000000000000110;
assign din[297] = 16'b0000000000010000;
assign din[298] = 16'b0000000001011010;
assign din[299] = 16'b0000000010111010;
assign din[300] = 16'b0000000011111001;
assign din[301] = 16'b0000000011110010;
assign din[302] = 16'b0000000010101001;
assign din[303] = 16'b0000000001001000;
assign din[304] = 16'b0000000000001000;
assign din[305] = 16'b0000000000001101;
assign din[306] = 16'b0000000001010100;
assign din[307] = 16'b0000000010110101;
assign din[308] = 16'b0000000011110111;
assign din[309] = 16'b0000000011110100;
assign din[310] = 16'b0000000010101111;
assign din[311] = 16'b0000000001001110;
assign din[312] = 16'b0000000000001011;
assign din[313] = 16'b0000000000001011;
assign din[314] = 16'b0000000001001110;
assign din[315] = 16'b0000000010101111;
assign din[316] = 16'b0000000011110100;
assign din[317] = 16'b0000000011110111;
assign din[318] = 16'b0000000010110101;
assign din[319] = 16'b0000000001010100;
assign din[320] = 16'b0000000000001101;
assign din[321] = 16'b0000000000001000;
assign din[322] = 16'b0000000001001000;
assign din[323] = 16'b0000000010101001;
assign din[324] = 16'b0000000011110010;
assign din[325] = 16'b0000000011111001;
assign din[326] = 16'b0000000010111010;
assign din[327] = 16'b0000000001011010;
assign din[328] = 16'b0000000000010000;
assign din[329] = 16'b0000000000000110;
assign din[330] = 16'b0000000001000011;
assign din[331] = 16'b0000000010100011;
assign din[332] = 16'b0000000011101111;
assign din[333] = 16'b0000000011111011;
assign din[334] = 16'b0000000011000000;
assign din[335] = 16'b0000000001100000;
assign din[336] = 16'b0000000000010011;
assign din[337] = 16'b0000000000000101;
assign din[338] = 16'b0000000000111101;
assign din[339] = 16'b0000000010011100;
assign din[340] = 16'b0000000011101011;
assign din[341] = 16'b0000000011111100;
assign din[342] = 16'b0000000011000101;
assign din[343] = 16'b0000000001100111;
assign din[344] = 16'b0000000000010111;
assign din[345] = 16'b0000000000000011;
assign din[346] = 16'b0000000000111000;
assign din[347] = 16'b0000000010010110;
assign din[348] = 16'b0000000011101000;
assign din[349] = 16'b0000000011111101;
assign din[350] = 16'b0000000011001011;
assign din[351] = 16'b0000000001101101;
assign din[352] = 16'b0000000000011010;
assign din[353] = 16'b0000000000000010;
assign din[354] = 16'b0000000000110011;
assign din[355] = 16'b0000000010010000;
assign din[356] = 16'b0000000011100100;
assign din[357] = 16'b0000000011111110;
assign din[358] = 16'b0000000011010000;
assign din[359] = 16'b0000000001110011;
assign din[360] = 16'b0000000000011110;
assign din[361] = 16'b0000000000000001;
assign din[362] = 16'b0000000000101110;
assign din[363] = 16'b0000000010001010;
assign din[364] = 16'b0000000011100000;
assign din[365] = 16'b0000000011111111;
assign din[366] = 16'b0000000011010101;
assign din[367] = 16'b0000000001111010;
assign din[368] = 16'b0000000000100010;
assign din[369] = 16'b0000000000000001;
assign din[370] = 16'b0000000000101001;
assign din[371] = 16'b0000000010000011;
assign din[372] = 16'b0000000011011011;
assign din[373] = 16'b0000000011111111;
assign din[374] = 16'b0000000011011001;
assign din[375] = 16'b0000000010000000;
assign din[376] = 16'b0000000000100111;
assign din[377] = 16'b0000000000000001;
assign din[378] = 16'b0000000000100101;
assign din[379] = 16'b0000000001111101;
assign din[380] = 16'b0000000011010111;
assign din[381] = 16'b0000000011111111;
assign din[382] = 16'b0000000011011110;
assign din[383] = 16'b0000000010000110;
assign din[384] = 16'b0000000000101011;
assign din[385] = 16'b0000000000000001;
assign din[386] = 16'b0000000000100000;
assign din[387] = 16'b0000000001110110;
assign din[388] = 16'b0000000011010010;
assign din[389] = 16'b0000000011111111;
assign din[390] = 16'b0000000011100010;
assign din[391] = 16'b0000000010001101;
assign din[392] = 16'b0000000000110000;
assign din[393] = 16'b0000000000000010;
assign din[394] = 16'b0000000000011100;
assign din[395] = 16'b0000000001110000;
assign din[396] = 16'b0000000011001101;
assign din[397] = 16'b0000000011111110;
assign din[398] = 16'b0000000011100110;
assign din[399] = 16'b0000000010010011;
assign din[400] = 16'b0000000000110101;
assign din[401] = 16'b0000000000000011;
assign din[402] = 16'b0000000000011000;
assign din[403] = 16'b0000000001101010;
assign din[404] = 16'b0000000011001000;
assign din[405] = 16'b0000000011111101;
assign din[406] = 16'b0000000011101001;
assign din[407] = 16'b0000000010011001;
assign din[408] = 16'b0000000000111011;
assign din[409] = 16'b0000000000000100;
assign din[410] = 16'b0000000000010101;
assign din[411] = 16'b0000000001100100;
assign din[412] = 16'b0000000011000011;
assign din[413] = 16'b0000000011111011;
assign din[414] = 16'b0000000011101101;
assign din[415] = 16'b0000000010100000;
assign din[416] = 16'b0000000001000000;
assign din[417] = 16'b0000000000000101;
assign din[418] = 16'b0000000000010001;
assign din[419] = 16'b0000000001011101;
assign din[420] = 16'b0000000010111101;
assign din[421] = 16'b0000000011111010;
assign din[422] = 16'b0000000011110000;
assign din[423] = 16'b0000000010100110;
assign din[424] = 16'b0000000001000110;
assign din[425] = 16'b0000000000000111;
assign din[426] = 16'b0000000000001110;
assign din[427] = 16'b0000000001010111;
assign din[428] = 16'b0000000010111000;
assign din[429] = 16'b0000000011111000;
assign din[430] = 16'b0000000011110011;
assign din[431] = 16'b0000000010101100;
assign din[432] = 16'b0000000001001011;
assign din[433] = 16'b0000000000001001;
assign din[434] = 16'b0000000000001100;
assign din[435] = 16'b0000000001010001;
assign din[436] = 16'b0000000010110010;
assign din[437] = 16'b0000000011110101;
assign din[438] = 16'b0000000011110101;
assign din[439] = 16'b0000000010110010;
assign din[440] = 16'b0000000001010001;
assign din[441] = 16'b0000000000001100;
assign din[442] = 16'b0000000000001001;
assign din[443] = 16'b0000000001001011;
assign din[444] = 16'b0000000010101100;
assign din[445] = 16'b0000000011110011;
assign din[446] = 16'b0000000011111000;
assign din[447] = 16'b0000000010111000;
assign din[448] = 16'b0000000001010111;
assign din[449] = 16'b0000000000001110;
assign din[450] = 16'b0000000000000111;
assign din[451] = 16'b0000000001000110;
assign din[452] = 16'b0000000010100110;
assign din[453] = 16'b0000000011110000;
assign din[454] = 16'b0000000011111010;
assign din[455] = 16'b0000000010111101;
assign din[456] = 16'b0000000001011101;
assign din[457] = 16'b0000000000010001;
assign din[458] = 16'b0000000000000101;
assign din[459] = 16'b0000000001000000;
assign din[460] = 16'b0000000010100000;
assign din[461] = 16'b0000000011101101;
assign din[462] = 16'b0000000011111011;
assign din[463] = 16'b0000000011000011;
assign din[464] = 16'b0000000001100100;
assign din[465] = 16'b0000000000010101;
assign din[466] = 16'b0000000000000100;
assign din[467] = 16'b0000000000111011;
assign din[468] = 16'b0000000010011001;
assign din[469] = 16'b0000000011101001;
assign din[470] = 16'b0000000011111101;
assign din[471] = 16'b0000000011001000;
assign din[472] = 16'b0000000001101010;
assign din[473] = 16'b0000000000011000;
assign din[474] = 16'b0000000000000011;
assign din[475] = 16'b0000000000110101;
assign din[476] = 16'b0000000010010011;
assign din[477] = 16'b0000000011100110;
assign din[478] = 16'b0000000011111110;
assign din[479] = 16'b0000000011001101;
assign din[480] = 16'b0000000001110000;
assign din[481] = 16'b0000000000011100;
assign din[482] = 16'b0000000000000010;
assign din[483] = 16'b0000000000110000;
assign din[484] = 16'b0000000010001101;
assign din[485] = 16'b0000000011100010;
assign din[486] = 16'b0000000011111111;
assign din[487] = 16'b0000000011010010;
assign din[488] = 16'b0000000001110110;
assign din[489] = 16'b0000000000100000;
assign din[490] = 16'b0000000000000001;
assign din[491] = 16'b0000000000101011;
assign din[492] = 16'b0000000010000110;
assign din[493] = 16'b0000000011011110;
assign din[494] = 16'b0000000011111111;
assign din[495] = 16'b0000000011010111;
assign din[496] = 16'b0000000001111101;
assign din[497] = 16'b0000000000100101;
assign din[498] = 16'b0000000000000001;
assign din[499] = 16'b0000000000100111;
assign din[500] = 16'b0000000010000000;
assign din[501] = 16'b0000000011011001;
assign din[502] = 16'b0000000011111111;
assign din[503] = 16'b0000000011011011;
assign din[504] = 16'b0000000010000011;
assign din[505] = 16'b0000000000101001;
assign din[506] = 16'b0000000000000001;
assign din[507] = 16'b0000000000100010;
assign din[508] = 16'b0000000001111010;
assign din[509] = 16'b0000000011010101;
assign din[510] = 16'b0000000011111111;
assign din[511] = 16'b0000000011100000;

assign din_out = din[add_rd];

endmodule