// whole note
// 20x30


module whole_note_rom (
    input logic clk,
    input logic [9:0] addr,
    output logic pixel_out
);


endmodule