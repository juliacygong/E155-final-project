// eighth note with upwards stem
// 20x30

module eighth_note_up_rom (
    input logic clk,
    input logic [9:0] addr,
    output logic pixel_out
);



endmodule