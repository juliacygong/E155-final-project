// Julia Gong
// 11/2/2025
// This file contains the lookup table for the twiddle factor values used in the FFT

module twiddleLUT(input logic [7:0] tw_add, // 8 bits good for 255
                  output logic [15:0] real_tw, // cos value
                  output logic [15:0] img_tw // sin value
                  );
				  

    // memory allocation buffer for real and imaginary twiddle factor values
    // 256 elements with 16 bit length
    logic [255:0][15:0] twiddle_cos;
    logic [255:0][15:0] twiddle_sin;

    // main LUT for twiddle addresses and values, where index [k] holds address
    // twiddle_cos = cos(2pi*k / 512)      twiddle_sin = sin(2pi*k / 512)

    assign twiddle_cos[0] = 16'h7FFF;      assign twiddle_sin[0] = 16'h0000; // cos: 1.000000, sin:0.000000
    assign twiddle_cos[1] = 16'h7FFD;      assign twiddle_sin[1] = 16'h0192; // cos: 0.999925, sin:0.012272
    assign twiddle_cos[2] = 16'h7FF5;      assign twiddle_sin[2] = 16'h0324; // cos: 0.999699, sin:0.024541
    assign twiddle_cos[3] = 16'h7FE9;      assign twiddle_sin[3] = 16'h04B6; // cos: 0.999322, sin:0.036807
    assign twiddle_cos[4] = 16'h7FD8;      assign twiddle_sin[4] = 16'h0648; // cos: 0.998795, sin:0.049068
    assign twiddle_cos[5] = 16'h7FC1;      assign twiddle_sin[5] = 16'h07D9; // cos: 0.998118, sin:0.061321
    assign twiddle_cos[6] = 16'h7FA6;      assign twiddle_sin[6] = 16'h096A; // cos: 0.997290, sin:0.073565
    assign twiddle_cos[7] = 16'h7F86;      assign twiddle_sin[7] = 16'h0AFB; // cos: 0.996313, sin:0.085797
    assign twiddle_cos[8] = 16'h7F61;      assign twiddle_sin[8] = 16'h0C8C; // cos: 0.995185, sin:0.098017
    assign twiddle_cos[9] = 16'h7F37;      assign twiddle_sin[9] = 16'h0E1C; // cos: 0.993907, sin:0.110222
    assign twiddle_cos[10] = 16'h7F09;      assign twiddle_sin[10] = 16'h0FAB; // cos: 0.992480, sin:0.122411
    assign twiddle_cos[11] = 16'h7ED5;      assign twiddle_sin[11] = 16'h113A; // cos: 0.990903, sin:0.134581
    assign twiddle_cos[12] = 16'h7E9C;      assign twiddle_sin[12] = 16'h12C8; // cos: 0.989177, sin:0.146730
    assign twiddle_cos[13] = 16'h7E5F;      assign twiddle_sin[13] = 16'h1455; // cos: 0.987301, sin:0.158858
    assign twiddle_cos[14] = 16'h7E1D;      assign twiddle_sin[14] = 16'h15E2; // cos: 0.985278, sin:0.170962
    assign twiddle_cos[15] = 16'h7DD5;      assign twiddle_sin[15] = 16'h176E; // cos: 0.983105, sin:0.183040
    assign twiddle_cos[16] = 16'h7D89;      assign twiddle_sin[16] = 16'h18F9; // cos: 0.980785, sin:0.195090
    assign twiddle_cos[17] = 16'h7D39;      assign twiddle_sin[17] = 16'h1A82; // cos: 0.978317, sin:0.207111
    assign twiddle_cos[18] = 16'h7CE3;      assign twiddle_sin[18] = 16'h1C0B; // cos: 0.975702, sin:0.219101
    assign twiddle_cos[19] = 16'h7C88;      assign twiddle_sin[19] = 16'h1D93; // cos: 0.972940, sin:0.231058
    assign twiddle_cos[20] = 16'h7C29;      assign twiddle_sin[20] = 16'h1F1A; // cos: 0.970031, sin:0.242980
    assign twiddle_cos[21] = 16'h7BC5;      assign twiddle_sin[21] = 16'h209F; // cos: 0.966976, sin:0.254866
    assign twiddle_cos[22] = 16'h7B5C;      assign twiddle_sin[22] = 16'h2223; // cos: 0.963776, sin:0.266713
    assign twiddle_cos[23] = 16'h7AEE;      assign twiddle_sin[23] = 16'h23A6; // cos: 0.960431, sin:0.278520
    assign twiddle_cos[24] = 16'h7A7C;      assign twiddle_sin[24] = 16'h2528; // cos: 0.956940, sin:0.290285
    assign twiddle_cos[25] = 16'h7A05;      assign twiddle_sin[25] = 16'h26A8; // cos: 0.953306, sin:0.302006
    assign twiddle_cos[26] = 16'h7989;      assign twiddle_sin[26] = 16'h2826; // cos: 0.949528, sin:0.313682
    assign twiddle_cos[27] = 16'h7909;      assign twiddle_sin[27] = 16'h29A3; // cos: 0.945607, sin:0.325310
    assign twiddle_cos[28] = 16'h7884;      assign twiddle_sin[28] = 16'h2B1F; // cos: 0.941544, sin:0.336890
    assign twiddle_cos[29] = 16'h77FA;      assign twiddle_sin[29] = 16'h2C99; // cos: 0.937339, sin:0.348419
    assign twiddle_cos[30] = 16'h776B;      assign twiddle_sin[30] = 16'h2E11; // cos: 0.932993, sin:0.359895
    assign twiddle_cos[31] = 16'h76D8;      assign twiddle_sin[31] = 16'h2F87; // cos: 0.928506, sin:0.371317
    assign twiddle_cos[32] = 16'h7641;      assign twiddle_sin[32] = 16'h30FB; // cos: 0.923880, sin:0.382683
    assign twiddle_cos[33] = 16'h75A5;      assign twiddle_sin[33] = 16'h326E; // cos: 0.919114, sin:0.393992
    assign twiddle_cos[34] = 16'h7504;      assign twiddle_sin[34] = 16'h33DF; // cos: 0.914210, sin:0.405241
    assign twiddle_cos[35] = 16'h745F;      assign twiddle_sin[35] = 16'h354D; // cos: 0.909168, sin:0.416430
    assign twiddle_cos[36] = 16'h73B5;      assign twiddle_sin[36] = 16'h36BA; // cos: 0.903989, sin:0.427555
    assign twiddle_cos[37] = 16'h7307;      assign twiddle_sin[37] = 16'h3824; // cos: 0.898674, sin:0.438616
    assign twiddle_cos[38] = 16'h7254;      assign twiddle_sin[38] = 16'h398C; // cos: 0.893224, sin:0.449611
    assign twiddle_cos[39] = 16'h719D;      assign twiddle_sin[39] = 16'h3AF2; // cos: 0.887640, sin:0.460539
    assign twiddle_cos[40] = 16'h70E2;      assign twiddle_sin[40] = 16'h3C56; // cos: 0.881921, sin:0.471397
    assign twiddle_cos[41] = 16'h7022;      assign twiddle_sin[41] = 16'h3DB8; // cos: 0.876070, sin:0.482184
    assign twiddle_cos[42] = 16'h6F5E;      assign twiddle_sin[42] = 16'h3F17; // cos: 0.870087, sin:0.492898
    assign twiddle_cos[43] = 16'h6E96;      assign twiddle_sin[43] = 16'h4073; // cos: 0.863973, sin:0.503538
    assign twiddle_cos[44] = 16'h6DC9;      assign twiddle_sin[44] = 16'h41CE; // cos: 0.857729, sin:0.514103
    assign twiddle_cos[45] = 16'h6CF8;      assign twiddle_sin[45] = 16'h4325; // cos: 0.851355, sin:0.524590
    assign twiddle_cos[46] = 16'h6C23;      assign twiddle_sin[46] = 16'h447A; // cos: 0.844854, sin:0.534998
    assign twiddle_cos[47] = 16'h6B4A;      assign twiddle_sin[47] = 16'h45CD; // cos: 0.838225, sin:0.545325
    assign twiddle_cos[48] = 16'h6A6D;      assign twiddle_sin[48] = 16'h471C; // cos: 0.831470, sin:0.555570
    assign twiddle_cos[49] = 16'h698B;      assign twiddle_sin[49] = 16'h4869; // cos: 0.824589, sin:0.565732
    assign twiddle_cos[50] = 16'h68A6;      assign twiddle_sin[50] = 16'h49B4; // cos: 0.817585, sin:0.575808
    assign twiddle_cos[51] = 16'h67BC;      assign twiddle_sin[51] = 16'h4AFB; // cos: 0.810457, sin:0.585798
    assign twiddle_cos[52] = 16'h66CF;      assign twiddle_sin[52] = 16'h4C3F; // cos: 0.803208, sin:0.595699
    assign twiddle_cos[53] = 16'h65DD;      assign twiddle_sin[53] = 16'h4D81; // cos: 0.795837, sin:0.605511
    assign twiddle_cos[54] = 16'h64E8;      assign twiddle_sin[54] = 16'h4EBF; // cos: 0.788346, sin:0.615232
    assign twiddle_cos[55] = 16'h63EE;      assign twiddle_sin[55] = 16'h4FFB; // cos: 0.780737, sin:0.624859
    assign twiddle_cos[56] = 16'h62F1;      assign twiddle_sin[56] = 16'h5133; // cos: 0.773010, sin:0.634393
    assign twiddle_cos[57] = 16'h61F0;      assign twiddle_sin[57] = 16'h5268; // cos: 0.765167, sin:0.643832
    assign twiddle_cos[58] = 16'h60EB;      assign twiddle_sin[58] = 16'h539B; // cos: 0.757209, sin:0.653173
    assign twiddle_cos[59] = 16'h5FE3;      assign twiddle_sin[59] = 16'h54C9; // cos: 0.749136, sin:0.662416
    assign twiddle_cos[60] = 16'h5ED7;      assign twiddle_sin[60] = 16'h55F5; // cos: 0.740951, sin:0.671559
    assign twiddle_cos[61] = 16'h5DC7;      assign twiddle_sin[61] = 16'h571D; // cos: 0.732654, sin:0.680601
    assign twiddle_cos[62] = 16'h5CB3;      assign twiddle_sin[62] = 16'h5842; // cos: 0.724247, sin:0.689541
    assign twiddle_cos[63] = 16'h5B9C;      assign twiddle_sin[63] = 16'h5964; // cos: 0.715731, sin:0.698376
    assign twiddle_cos[64] = 16'h5A82;      assign twiddle_sin[64] = 16'h5A82; // cos: 0.707107, sin:0.707107
    assign twiddle_cos[65] = 16'h5964;      assign twiddle_sin[65] = 16'h5B9C; // cos: 0.698376, sin:0.715731
    assign twiddle_cos[66] = 16'h5842;      assign twiddle_sin[66] = 16'h5CB3; // cos: 0.689541, sin:0.724247
    assign twiddle_cos[67] = 16'h571D;      assign twiddle_sin[67] = 16'h5DC7; // cos: 0.680601, sin:0.732654
    assign twiddle_cos[68] = 16'h55F5;      assign twiddle_sin[68] = 16'h5ED7; // cos: 0.671559, sin:0.740951
    assign twiddle_cos[69] = 16'h54C9;      assign twiddle_sin[69] = 16'h5FE3; // cos: 0.662416, sin:0.749136
    assign twiddle_cos[70] = 16'h539B;      assign twiddle_sin[70] = 16'h60EB; // cos: 0.653173, sin:0.757209
    assign twiddle_cos[71] = 16'h5268;      assign twiddle_sin[71] = 16'h61F0; // cos: 0.643832, sin:0.765167
    assign twiddle_cos[72] = 16'h5133;      assign twiddle_sin[72] = 16'h62F1; // cos: 0.634393, sin:0.773010
    assign twiddle_cos[73] = 16'h4FFB;      assign twiddle_sin[73] = 16'h63EE; // cos: 0.624859, sin:0.780737
    assign twiddle_cos[74] = 16'h4EBF;      assign twiddle_sin[74] = 16'h64E8; // cos: 0.615232, sin:0.788346
    assign twiddle_cos[75] = 16'h4D81;      assign twiddle_sin[75] = 16'h65DD; // cos: 0.605511, sin:0.795837
    assign twiddle_cos[76] = 16'h4C3F;      assign twiddle_sin[76] = 16'h66CF; // cos: 0.595699, sin:0.803208
    assign twiddle_cos[77] = 16'h4AFB;      assign twiddle_sin[77] = 16'h67BC; // cos: 0.585798, sin:0.810457
    assign twiddle_cos[78] = 16'h49B4;      assign twiddle_sin[78] = 16'h68A6; // cos: 0.575808, sin:0.817585
    assign twiddle_cos[79] = 16'h4869;      assign twiddle_sin[79] = 16'h698B; // cos: 0.565732, sin:0.824589
    assign twiddle_cos[80] = 16'h471C;      assign twiddle_sin[80] = 16'h6A6D; // cos: 0.555570, sin:0.831470
    assign twiddle_cos[81] = 16'h45CD;      assign twiddle_sin[81] = 16'h6B4A; // cos: 0.545325, sin:0.838225
    assign twiddle_cos[82] = 16'h447A;      assign twiddle_sin[82] = 16'h6C23; // cos: 0.534998, sin:0.844854
    assign twiddle_cos[83] = 16'h4325;      assign twiddle_sin[83] = 16'h6CF8; // cos: 0.524590, sin:0.851355
    assign twiddle_cos[84] = 16'h41CE;      assign twiddle_sin[84] = 16'h6DC9; // cos: 0.514103, sin:0.857729
    assign twiddle_cos[85] = 16'h4073;      assign twiddle_sin[85] = 16'h6E96; // cos: 0.503538, sin:0.863973
    assign twiddle_cos[86] = 16'h3F17;      assign twiddle_sin[86] = 16'h6F5E; // cos: 0.492898, sin:0.870087
    assign twiddle_cos[87] = 16'h3DB8;      assign twiddle_sin[87] = 16'h7022; // cos: 0.482184, sin:0.876070
    assign twiddle_cos[88] = 16'h3C56;      assign twiddle_sin[88] = 16'h70E2; // cos: 0.471397, sin:0.881921
    assign twiddle_cos[89] = 16'h3AF2;      assign twiddle_sin[89] = 16'h719D; // cos: 0.460539, sin:0.887640
    assign twiddle_cos[90] = 16'h398C;      assign twiddle_sin[90] = 16'h7254; // cos: 0.449611, sin:0.893224
    assign twiddle_cos[91] = 16'h3824;      assign twiddle_sin[91] = 16'h7307; // cos: 0.438616, sin:0.898674
    assign twiddle_cos[92] = 16'h36BA;      assign twiddle_sin[92] = 16'h73B5; // cos: 0.427555, sin:0.903989
    assign twiddle_cos[93] = 16'h354D;      assign twiddle_sin[93] = 16'h745F; // cos: 0.416430, sin:0.909168
    assign twiddle_cos[94] = 16'h33DF;      assign twiddle_sin[94] = 16'h7504; // cos: 0.405241, sin:0.914210
    assign twiddle_cos[95] = 16'h326E;      assign twiddle_sin[95] = 16'h75A5; // cos: 0.393992, sin:0.919114
    assign twiddle_cos[96] = 16'h30FB;      assign twiddle_sin[96] = 16'h7641; // cos: 0.382683, sin:0.923880
    assign twiddle_cos[97] = 16'h2F87;      assign twiddle_sin[97] = 16'h76D8; // cos: 0.371317, sin:0.928506
    assign twiddle_cos[98] = 16'h2E11;      assign twiddle_sin[98] = 16'h776B; // cos: 0.359895, sin:0.932993
    assign twiddle_cos[99] = 16'h2C99;      assign twiddle_sin[99] = 16'h77FA; // cos: 0.348419, sin:0.937339
    assign twiddle_cos[100] = 16'h2B1F;      assign twiddle_sin[100] = 16'h7884; // cos: 0.336890, sin:0.941544
    assign twiddle_cos[101] = 16'h29A3;      assign twiddle_sin[101] = 16'h7909; // cos: 0.325310, sin:0.945607
    assign twiddle_cos[102] = 16'h2826;      assign twiddle_sin[102] = 16'h7989; // cos: 0.313682, sin:0.949528
    assign twiddle_cos[103] = 16'h26A8;      assign twiddle_sin[103] = 16'h7A05; // cos: 0.302006, sin:0.953306
    assign twiddle_cos[104] = 16'h2528;      assign twiddle_sin[104] = 16'h7A7C; // cos: 0.290285, sin:0.956940
    assign twiddle_cos[105] = 16'h23A6;      assign twiddle_sin[105] = 16'h7AEE; // cos: 0.278520, sin:0.960431
    assign twiddle_cos[106] = 16'h2223;      assign twiddle_sin[106] = 16'h7B5C; // cos: 0.266713, sin:0.963776
    assign twiddle_cos[107] = 16'h209F;      assign twiddle_sin[107] = 16'h7BC5; // cos: 0.254866, sin:0.966976
    assign twiddle_cos[108] = 16'h1F1A;      assign twiddle_sin[108] = 16'h7C29; // cos: 0.242980, sin:0.970031
    assign twiddle_cos[109] = 16'h1D93;      assign twiddle_sin[109] = 16'h7C88; // cos: 0.231058, sin:0.972940
    assign twiddle_cos[110] = 16'h1C0B;      assign twiddle_sin[110] = 16'h7CE3; // cos: 0.219101, sin:0.975702
    assign twiddle_cos[111] = 16'h1A82;      assign twiddle_sin[111] = 16'h7D39; // cos: 0.207111, sin:0.978317
    assign twiddle_cos[112] = 16'h18F9;      assign twiddle_sin[112] = 16'h7D89; // cos: 0.195090, sin:0.980785
    assign twiddle_cos[113] = 16'h176E;      assign twiddle_sin[113] = 16'h7DD5; // cos: 0.183040, sin:0.983105
    assign twiddle_cos[114] = 16'h15E2;      assign twiddle_sin[114] = 16'h7E1D; // cos: 0.170962, sin:0.985278
    assign twiddle_cos[115] = 16'h1455;      assign twiddle_sin[115] = 16'h7E5F; // cos: 0.158858, sin:0.987301
    assign twiddle_cos[116] = 16'h12C8;      assign twiddle_sin[116] = 16'h7E9C; // cos: 0.146730, sin:0.989177
    assign twiddle_cos[117] = 16'h113A;      assign twiddle_sin[117] = 16'h7ED5; // cos: 0.134581, sin:0.990903
    assign twiddle_cos[118] = 16'h0FAB;      assign twiddle_sin[118] = 16'h7F09; // cos: 0.122411, sin:0.992480
    assign twiddle_cos[119] = 16'h0E1C;      assign twiddle_sin[119] = 16'h7F37; // cos: 0.110222, sin:0.993907
    assign twiddle_cos[120] = 16'h0C8C;      assign twiddle_sin[120] = 16'h7F61; // cos: 0.098017, sin:0.995185
    assign twiddle_cos[121] = 16'h0AFB;      assign twiddle_sin[121] = 16'h7F86; // cos: 0.085797, sin:0.996313
    assign twiddle_cos[122] = 16'h096A;      assign twiddle_sin[122] = 16'h7FA6; // cos: 0.073565, sin:0.997290
    assign twiddle_cos[123] = 16'h07D9;      assign twiddle_sin[123] = 16'h7FC1; // cos: 0.061321, sin:0.998118
    assign twiddle_cos[124] = 16'h0648;      assign twiddle_sin[124] = 16'h7FD8; // cos: 0.049068, sin:0.998795
    assign twiddle_cos[125] = 16'h04B6;      assign twiddle_sin[125] = 16'h7FE9; // cos: 0.036807, sin:0.999322
    assign twiddle_cos[126] = 16'h0324;      assign twiddle_sin[126] = 16'h7FF5; // cos: 0.024541, sin:0.999699
    assign twiddle_cos[127] = 16'h0192;      assign twiddle_sin[127] = 16'h7FFD; // cos: 0.012272, sin:0.999925
    assign twiddle_cos[128] = 16'h0000;      assign twiddle_sin[128] = 16'h7FFF; // cos: 0.000000, sin:1.000000
    assign twiddle_cos[129] = 16'hFE6E;      assign twiddle_sin[129] = 16'h7FFD; // cos: -0.012272, sin:0.999925
    assign twiddle_cos[130] = 16'hFCDC;      assign twiddle_sin[130] = 16'h7FF5; // cos: -0.024541, sin:0.999699
    assign twiddle_cos[131] = 16'hFB4A;      assign twiddle_sin[131] = 16'h7FE9; // cos: -0.036807, sin:0.999322
    assign twiddle_cos[132] = 16'hF9B8;      assign twiddle_sin[132] = 16'h7FD8; // cos: -0.049068, sin:0.998795
    assign twiddle_cos[133] = 16'hF827;      assign twiddle_sin[133] = 16'h7FC1; // cos: -0.061321, sin:0.998118
    assign twiddle_cos[134] = 16'hF696;      assign twiddle_sin[134] = 16'h7FA6; // cos: -0.073565, sin:0.997290
    assign twiddle_cos[135] = 16'hF505;      assign twiddle_sin[135] = 16'h7F86; // cos: -0.085797, sin:0.996313
    assign twiddle_cos[136] = 16'hF374;      assign twiddle_sin[136] = 16'h7F61; // cos: -0.098017, sin:0.995185
    assign twiddle_cos[137] = 16'hF1E4;      assign twiddle_sin[137] = 16'h7F37; // cos: -0.110222, sin:0.993907
    assign twiddle_cos[138] = 16'hF055;      assign twiddle_sin[138] = 16'h7F09; // cos: -0.122411, sin:0.992480
    assign twiddle_cos[139] = 16'hEEC6;      assign twiddle_sin[139] = 16'h7ED5; // cos: -0.134581, sin:0.990903
    assign twiddle_cos[140] = 16'hED38;      assign twiddle_sin[140] = 16'h7E9C; // cos: -0.146730, sin:0.989177
    assign twiddle_cos[141] = 16'hEBAB;      assign twiddle_sin[141] = 16'h7E5F; // cos: -0.158858, sin:0.987301
    assign twiddle_cos[142] = 16'hEA1E;      assign twiddle_sin[142] = 16'h7E1D; // cos: -0.170962, sin:0.985278
    assign twiddle_cos[143] = 16'hE892;      assign twiddle_sin[143] = 16'h7DD5; // cos: -0.183040, sin:0.983105
    assign twiddle_cos[144] = 16'hE707;      assign twiddle_sin[144] = 16'h7D89; // cos: -0.195090, sin:0.980785
    assign twiddle_cos[145] = 16'hE57E;      assign twiddle_sin[145] = 16'h7D39; // cos: -0.207111, sin:0.978317
    assign twiddle_cos[146] = 16'hE3F5;      assign twiddle_sin[146] = 16'h7CE3; // cos: -0.219101, sin:0.975702
    assign twiddle_cos[147] = 16'hE26D;      assign twiddle_sin[147] = 16'h7C88; // cos: -0.231058, sin:0.972940
    assign twiddle_cos[148] = 16'hE0E6;      assign twiddle_sin[148] = 16'h7C29; // cos: -0.242980, sin:0.970031
    assign twiddle_cos[149] = 16'hDF61;      assign twiddle_sin[149] = 16'h7BC5; // cos: -0.254866, sin:0.966976
    assign twiddle_cos[150] = 16'hDDDD;      assign twiddle_sin[150] = 16'h7B5C; // cos: -0.266713, sin:0.963776
    assign twiddle_cos[151] = 16'hDC5A;      assign twiddle_sin[151] = 16'h7AEE; // cos: -0.278520, sin:0.960431
    assign twiddle_cos[152] = 16'hDAD8;      assign twiddle_sin[152] = 16'h7A7C; // cos: -0.290285, sin:0.956940
    assign twiddle_cos[153] = 16'hD958;      assign twiddle_sin[153] = 16'h7A05; // cos: -0.302006, sin:0.953306
    assign twiddle_cos[154] = 16'hD7DA;      assign twiddle_sin[154] = 16'h7989; // cos: -0.313682, sin:0.949528
    assign twiddle_cos[155] = 16'hD65D;      assign twiddle_sin[155] = 16'h7909; // cos: -0.325310, sin:0.945607
    assign twiddle_cos[156] = 16'hD4E1;      assign twiddle_sin[156] = 16'h7884; // cos: -0.336890, sin:0.941544
    assign twiddle_cos[157] = 16'hD367;      assign twiddle_sin[157] = 16'h77FA; // cos: -0.348419, sin:0.937339
    assign twiddle_cos[158] = 16'hD1EF;      assign twiddle_sin[158] = 16'h776B; // cos: -0.359895, sin:0.932993
    assign twiddle_cos[159] = 16'hD079;      assign twiddle_sin[159] = 16'h76D8; // cos: -0.371317, sin:0.928506
    assign twiddle_cos[160] = 16'hCF05;      assign twiddle_sin[160] = 16'h7641; // cos: -0.382683, sin:0.923880
    assign twiddle_cos[161] = 16'hCD92;      assign twiddle_sin[161] = 16'h75A5; // cos: -0.393992, sin:0.919114
    assign twiddle_cos[162] = 16'hCC21;      assign twiddle_sin[162] = 16'h7504; // cos: -0.405241, sin:0.914210
    assign twiddle_cos[163] = 16'hCAB3;      assign twiddle_sin[163] = 16'h745F; // cos: -0.416430, sin:0.909168
    assign twiddle_cos[164] = 16'hC946;      assign twiddle_sin[164] = 16'h73B5; // cos: -0.427555, sin:0.903989
    assign twiddle_cos[165] = 16'hC7DC;      assign twiddle_sin[165] = 16'h7307; // cos: -0.438616, sin:0.898674
    assign twiddle_cos[166] = 16'hC674;      assign twiddle_sin[166] = 16'h7254; // cos: -0.449611, sin:0.893224
    assign twiddle_cos[167] = 16'hC50E;      assign twiddle_sin[167] = 16'h719D; // cos: -0.460539, sin:0.887640
    assign twiddle_cos[168] = 16'hC3AA;      assign twiddle_sin[168] = 16'h70E2; // cos: -0.471397, sin:0.881921
    assign twiddle_cos[169] = 16'hC248;      assign twiddle_sin[169] = 16'h7022; // cos: -0.482184, sin:0.876070
    assign twiddle_cos[170] = 16'hC0E9;      assign twiddle_sin[170] = 16'h6F5E; // cos: -0.492898, sin:0.870087
    assign twiddle_cos[171] = 16'hBF8D;      assign twiddle_sin[171] = 16'h6E96; // cos: -0.503538, sin:0.863973
    assign twiddle_cos[172] = 16'hBE32;      assign twiddle_sin[172] = 16'h6DC9; // cos: -0.514103, sin:0.857729
    assign twiddle_cos[173] = 16'hBCDB;      assign twiddle_sin[173] = 16'h6CF8; // cos: -0.524590, sin:0.851355
    assign twiddle_cos[174] = 16'hBB86;      assign twiddle_sin[174] = 16'h6C23; // cos: -0.534998, sin:0.844854
    assign twiddle_cos[175] = 16'hBA33;      assign twiddle_sin[175] = 16'h6B4A; // cos: -0.545325, sin:0.838225
    assign twiddle_cos[176] = 16'hB8E4;      assign twiddle_sin[176] = 16'h6A6D; // cos: -0.555570, sin:0.831470
    assign twiddle_cos[177] = 16'hB797;      assign twiddle_sin[177] = 16'h698B; // cos: -0.565732, sin:0.824589
    assign twiddle_cos[178] = 16'hB64C;      assign twiddle_sin[178] = 16'h68A6; // cos: -0.575808, sin:0.817585
    assign twiddle_cos[179] = 16'hB505;      assign twiddle_sin[179] = 16'h67BC; // cos: -0.585798, sin:0.810457
    assign twiddle_cos[180] = 16'hB3C1;      assign twiddle_sin[180] = 16'h66CF; // cos: -0.595699, sin:0.803208
    assign twiddle_cos[181] = 16'hB27F;      assign twiddle_sin[181] = 16'h65DD; // cos: -0.605511, sin:0.795837
    assign twiddle_cos[182] = 16'hB141;      assign twiddle_sin[182] = 16'h64E8; // cos: -0.615232, sin:0.788346
    assign twiddle_cos[183] = 16'hB005;      assign twiddle_sin[183] = 16'h63EE; // cos: -0.624859, sin:0.780737
    assign twiddle_cos[184] = 16'hAECD;      assign twiddle_sin[184] = 16'h62F1; // cos: -0.634393, sin:0.773010
    assign twiddle_cos[185] = 16'hAD98;      assign twiddle_sin[185] = 16'h61F0; // cos: -0.643832, sin:0.765167
    assign twiddle_cos[186] = 16'hAC65;      assign twiddle_sin[186] = 16'h60EB; // cos: -0.653173, sin:0.757209
    assign twiddle_cos[187] = 16'hAB37;      assign twiddle_sin[187] = 16'h5FE3; // cos: -0.662416, sin:0.749136
    assign twiddle_cos[188] = 16'hAA0B;      assign twiddle_sin[188] = 16'h5ED7; // cos: -0.671559, sin:0.740951
    assign twiddle_cos[189] = 16'hA8E3;      assign twiddle_sin[189] = 16'h5DC7; // cos: -0.680601, sin:0.732654
    assign twiddle_cos[190] = 16'hA7BE;      assign twiddle_sin[190] = 16'h5CB3; // cos: -0.689541, sin:0.724247
    assign twiddle_cos[191] = 16'hA69C;      assign twiddle_sin[191] = 16'h5B9C; // cos: -0.698376, sin:0.715731
    assign twiddle_cos[192] = 16'hA57E;      assign twiddle_sin[192] = 16'h5A82; // cos: -0.707107, sin:0.707107
    assign twiddle_cos[193] = 16'hA464;      assign twiddle_sin[193] = 16'h5964; // cos: -0.715731, sin:0.698376
    assign twiddle_cos[194] = 16'hA34D;      assign twiddle_sin[194] = 16'h5842; // cos: -0.724247, sin:0.689541
    assign twiddle_cos[195] = 16'hA239;      assign twiddle_sin[195] = 16'h571D; // cos: -0.732654, sin:0.680601
    assign twiddle_cos[196] = 16'hA129;      assign twiddle_sin[196] = 16'h55F5; // cos: -0.740951, sin:0.671559
    assign twiddle_cos[197] = 16'hA01D;      assign twiddle_sin[197] = 16'h54C9; // cos: -0.749136, sin:0.662416
    assign twiddle_cos[198] = 16'h9F15;      assign twiddle_sin[198] = 16'h539B; // cos: -0.757209, sin:0.653173
    assign twiddle_cos[199] = 16'h9E10;      assign twiddle_sin[199] = 16'h5268; // cos: -0.765167, sin:0.643832
    assign twiddle_cos[200] = 16'h9D0F;      assign twiddle_sin[200] = 16'h5133; // cos: -0.773010, sin:0.634393
    assign twiddle_cos[201] = 16'h9C12;      assign twiddle_sin[201] = 16'h4FFB; // cos: -0.780737, sin:0.624859
    assign twiddle_cos[202] = 16'h9B18;      assign twiddle_sin[202] = 16'h4EBF; // cos: -0.788346, sin:0.615232
    assign twiddle_cos[203] = 16'h9A23;      assign twiddle_sin[203] = 16'h4D81; // cos: -0.795837, sin:0.605511
    assign twiddle_cos[204] = 16'h9931;      assign twiddle_sin[204] = 16'h4C3F; // cos: -0.803208, sin:0.595699
    assign twiddle_cos[205] = 16'h9844;      assign twiddle_sin[205] = 16'h4AFB; // cos: -0.810457, sin:0.585798
    assign twiddle_cos[206] = 16'h975A;      assign twiddle_sin[206] = 16'h49B4; // cos: -0.817585, sin:0.575808
    assign twiddle_cos[207] = 16'h9675;      assign twiddle_sin[207] = 16'h4869; // cos: -0.824589, sin:0.565732
    assign twiddle_cos[208] = 16'h9593;      assign twiddle_sin[208] = 16'h471C; // cos: -0.831470, sin:0.555570
    assign twiddle_cos[209] = 16'h94B6;      assign twiddle_sin[209] = 16'h45CD; // cos: -0.838225, sin:0.545325
    assign twiddle_cos[210] = 16'h93DD;      assign twiddle_sin[210] = 16'h447A; // cos: -0.844854, sin:0.534998
    assign twiddle_cos[211] = 16'h9308;      assign twiddle_sin[211] = 16'h4325; // cos: -0.851355, sin:0.524590
    assign twiddle_cos[212] = 16'h9237;      assign twiddle_sin[212] = 16'h41CE; // cos: -0.857729, sin:0.514103
    assign twiddle_cos[213] = 16'h916A;      assign twiddle_sin[213] = 16'h4073; // cos: -0.863973, sin:0.503538
    assign twiddle_cos[214] = 16'h90A2;      assign twiddle_sin[214] = 16'h3F17; // cos: -0.870087, sin:0.492898
    assign twiddle_cos[215] = 16'h8FDE;      assign twiddle_sin[215] = 16'h3DB8; // cos: -0.876070, sin:0.482184
    assign twiddle_cos[216] = 16'h8F1E;      assign twiddle_sin[216] = 16'h3C56; // cos: -0.881921, sin:0.471397
    assign twiddle_cos[217] = 16'h8E63;      assign twiddle_sin[217] = 16'h3AF2; // cos: -0.887640, sin:0.460539
    assign twiddle_cos[218] = 16'h8DAC;      assign twiddle_sin[218] = 16'h398C; // cos: -0.893224, sin:0.449611
    assign twiddle_cos[219] = 16'h8CF9;      assign twiddle_sin[219] = 16'h3824; // cos: -0.898674, sin:0.438616
    assign twiddle_cos[220] = 16'h8C4B;      assign twiddle_sin[220] = 16'h36BA; // cos: -0.903989, sin:0.427555
    assign twiddle_cos[221] = 16'h8BA1;      assign twiddle_sin[221] = 16'h354D; // cos: -0.909168, sin:0.416430
    assign twiddle_cos[222] = 16'h8AFC;      assign twiddle_sin[222] = 16'h33DF; // cos: -0.914210, sin:0.405241
    assign twiddle_cos[223] = 16'h8A5B;      assign twiddle_sin[223] = 16'h326E; // cos: -0.919114, sin:0.393992
    assign twiddle_cos[224] = 16'h89BF;      assign twiddle_sin[224] = 16'h30FB; // cos: -0.923880, sin:0.382683
    assign twiddle_cos[225] = 16'h8928;      assign twiddle_sin[225] = 16'h2F87; // cos: -0.928506, sin:0.371317
    assign twiddle_cos[226] = 16'h8895;      assign twiddle_sin[226] = 16'h2E11; // cos: -0.932993, sin:0.359895
    assign twiddle_cos[227] = 16'h8806;      assign twiddle_sin[227] = 16'h2C99; // cos: -0.937339, sin:0.348419
    assign twiddle_cos[228] = 16'h877C;      assign twiddle_sin[228] = 16'h2B1F; // cos: -0.941544, sin:0.336890
    assign twiddle_cos[229] = 16'h86F7;      assign twiddle_sin[229] = 16'h29A3; // cos: -0.945607, sin:0.325310
    assign twiddle_cos[230] = 16'h8677;      assign twiddle_sin[230] = 16'h2826; // cos: -0.949528, sin:0.313682
    assign twiddle_cos[231] = 16'h85FB;      assign twiddle_sin[231] = 16'h26A8; // cos: -0.953306, sin:0.302006
    assign twiddle_cos[232] = 16'h8584;      assign twiddle_sin[232] = 16'h2528; // cos: -0.956940, sin:0.290285
    assign twiddle_cos[233] = 16'h8512;      assign twiddle_sin[233] = 16'h23A6; // cos: -0.960431, sin:0.278520
    assign twiddle_cos[234] = 16'h84A4;      assign twiddle_sin[234] = 16'h2223; // cos: -0.963776, sin:0.266713
    assign twiddle_cos[235] = 16'h843B;      assign twiddle_sin[235] = 16'h209F; // cos: -0.966976, sin:0.254866
    assign twiddle_cos[236] = 16'h83D7;      assign twiddle_sin[236] = 16'h1F1A; // cos: -0.970031, sin:0.242980
    assign twiddle_cos[237] = 16'h8378;      assign twiddle_sin[237] = 16'h1D93; // cos: -0.972940, sin:0.231058
    assign twiddle_cos[238] = 16'h831D;      assign twiddle_sin[238] = 16'h1C0B; // cos: -0.975702, sin:0.219101
    assign twiddle_cos[239] = 16'h82C7;      assign twiddle_sin[239] = 16'h1A82; // cos: -0.978317, sin:0.207111
    assign twiddle_cos[240] = 16'h8277;      assign twiddle_sin[240] = 16'h18F9; // cos: -0.980785, sin:0.195090
    assign twiddle_cos[241] = 16'h822B;      assign twiddle_sin[241] = 16'h176E; // cos: -0.983105, sin:0.183040
    assign twiddle_cos[242] = 16'h81E3;      assign twiddle_sin[242] = 16'h15E2; // cos: -0.985278, sin:0.170962
    assign twiddle_cos[243] = 16'h81A1;      assign twiddle_sin[243] = 16'h1455; // cos: -0.987301, sin:0.158858
    assign twiddle_cos[244] = 16'h8164;      assign twiddle_sin[244] = 16'h12C8; // cos: -0.989177, sin:0.146730
    assign twiddle_cos[245] = 16'h812B;      assign twiddle_sin[245] = 16'h113A; // cos: -0.990903, sin:0.134581
    assign twiddle_cos[246] = 16'h80F7;      assign twiddle_sin[246] = 16'h0FAB; // cos: -0.992480, sin:0.122411
    assign twiddle_cos[247] = 16'h80C9;      assign twiddle_sin[247] = 16'h0E1C; // cos: -0.993907, sin:0.110222
    assign twiddle_cos[248] = 16'h809F;      assign twiddle_sin[248] = 16'h0C8C; // cos: -0.995185, sin:0.098017
    assign twiddle_cos[249] = 16'h807A;      assign twiddle_sin[249] = 16'h0AFB; // cos: -0.996313, sin:0.085797
    assign twiddle_cos[250] = 16'h805A;      assign twiddle_sin[250] = 16'h096A; // cos: -0.997290, sin:0.073565
    assign twiddle_cos[251] = 16'h803F;      assign twiddle_sin[251] = 16'h07D9; // cos: -0.998118, sin:0.061321
    assign twiddle_cos[252] = 16'h8028;      assign twiddle_sin[252] = 16'h0648; // cos: -0.998795, sin:0.049068
    assign twiddle_cos[253] = 16'h8017;      assign twiddle_sin[253] = 16'h04B6; // cos: -0.999322, sin:0.036807
    assign twiddle_cos[254] = 16'h800B;      assign twiddle_sin[254] = 16'h0324; // cos: -0.999699, sin:0.024541
    assign twiddle_cos[255] = 16'h8003;      assign twiddle_sin[255] = 16'h0192; // cos: -0.999925, sin:0.012272
	
	assign real_tw = twiddle_cos[tw_add];
	assign img_tw = -twiddle_sin[tw_add];

    endmodule